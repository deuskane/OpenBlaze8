library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity soft/identity is
  port (
    clk_i    : in std_logic;
    addr_i   : in std_logic_vector(9 downto 0);
    data_o   : out std_logic_vector(17 downto 0)
  );
end soft/identity ;

architecture behavioral of soft/identity is
begin
  read : process(clk_i)
  begin
    if(clk_i'event and clk_i = '1') then
      case to_integer(unsigned(addr_i)) is
        when 0 => data_o <= "000100000000000000";
        when 1 => data_o <= "101100000000000100";
        when 2 => data_o <= "110100000000000000";
        when 3 => data_o <= "000000000000000000";
        when 4 => data_o <= "000000000000000000";
        when 5 => data_o <= "000000000000000000";
        when 6 => data_o <= "000000000000000000";
        when 7 => data_o <= "000000000000000000";
        when 8 => data_o <= "000000000000000000";
        when 9 => data_o <= "000000000000000000";
        when 10 => data_o <= "000000000000000000";
        when 11 => data_o <= "000000000000000000";
        when 12 => data_o <= "000000000000000000";
        when 13 => data_o <= "000000000000000000";
        when 14 => data_o <= "000000000000000000";
        when 15 => data_o <= "000000000000000000";
        when 16 => data_o <= "000000000000000000";
        when 17 => data_o <= "000000000000000000";
        when 18 => data_o <= "000000000000000000";
        when 19 => data_o <= "000000000000000000";
        when 20 => data_o <= "000000000000000000";
        when 21 => data_o <= "000000000000000000";
        when 22 => data_o <= "000000000000000000";
        when 23 => data_o <= "000000000000000000";
        when 24 => data_o <= "000000000000000000";
        when 25 => data_o <= "000000000000000000";
        when 26 => data_o <= "000000000000000000";
        when 27 => data_o <= "000000000000000000";
        when 28 => data_o <= "000000000000000000";
        when 29 => data_o <= "000000000000000000";
        when 30 => data_o <= "000000000000000000";
        when 31 => data_o <= "000000000000000000";
        when 32 => data_o <= "000000000000000000";
        when 33 => data_o <= "000000000000000000";
        when 34 => data_o <= "000000000000000000";
        when 35 => data_o <= "000000000000000000";
        when 36 => data_o <= "000000000000000000";
        when 37 => data_o <= "000000000000000000";
        when 38 => data_o <= "000000000000000000";
        when 39 => data_o <= "000000000000000000";
        when 40 => data_o <= "000000000000000000";
        when 41 => data_o <= "000000000000000000";
        when 42 => data_o <= "000000000000000000";
        when 43 => data_o <= "000000000000000000";
        when 44 => data_o <= "000000000000000000";
        when 45 => data_o <= "000000000000000000";
        when 46 => data_o <= "000000000000000000";
        when 47 => data_o <= "000000000000000000";
        when 48 => data_o <= "000000000000000000";
        when 49 => data_o <= "000000000000000000";
        when 50 => data_o <= "000000000000000000";
        when 51 => data_o <= "000000000000000000";
        when 52 => data_o <= "000000000000000000";
        when 53 => data_o <= "000000000000000000";
        when 54 => data_o <= "000000000000000000";
        when 55 => data_o <= "000000000000000000";
        when 56 => data_o <= "000000000000000000";
        when 57 => data_o <= "000000000000000000";
        when 58 => data_o <= "000000000000000000";
        when 59 => data_o <= "000000000000000000";
        when 60 => data_o <= "000000000000000000";
        when 61 => data_o <= "000000000000000000";
        when 62 => data_o <= "000000000000000000";
        when 63 => data_o <= "000000000000000000";
        when 64 => data_o <= "000000000000000000";
        when 65 => data_o <= "000000000000000000";
        when 66 => data_o <= "000000000000000000";
        when 67 => data_o <= "000000000000000000";
        when 68 => data_o <= "000000000000000000";
        when 69 => data_o <= "000000000000000000";
        when 70 => data_o <= "000000000000000000";
        when 71 => data_o <= "000000000000000000";
        when 72 => data_o <= "000000000000000000";
        when 73 => data_o <= "000000000000000000";
        when 74 => data_o <= "000000000000000000";
        when 75 => data_o <= "000000000000000000";
        when 76 => data_o <= "000000000000000000";
        when 77 => data_o <= "000000000000000000";
        when 78 => data_o <= "000000000000000000";
        when 79 => data_o <= "000000000000000000";
        when 80 => data_o <= "000000000000000000";
        when 81 => data_o <= "000000000000000000";
        when 82 => data_o <= "000000000000000000";
        when 83 => data_o <= "000000000000000000";
        when 84 => data_o <= "000000000000000000";
        when 85 => data_o <= "000000000000000000";
        when 86 => data_o <= "000000000000000000";
        when 87 => data_o <= "000000000000000000";
        when 88 => data_o <= "000000000000000000";
        when 89 => data_o <= "000000000000000000";
        when 90 => data_o <= "000000000000000000";
        when 91 => data_o <= "000000000000000000";
        when 92 => data_o <= "000000000000000000";
        when 93 => data_o <= "000000000000000000";
        when 94 => data_o <= "000000000000000000";
        when 95 => data_o <= "000000000000000000";
        when 96 => data_o <= "000000000000000000";
        when 97 => data_o <= "000000000000000000";
        when 98 => data_o <= "000000000000000000";
        when 99 => data_o <= "000000000000000000";
        when 100 => data_o <= "000000000000000000";
        when 101 => data_o <= "000000000000000000";
        when 102 => data_o <= "000000000000000000";
        when 103 => data_o <= "000000000000000000";
        when 104 => data_o <= "000000000000000000";
        when 105 => data_o <= "000000000000000000";
        when 106 => data_o <= "000000000000000000";
        when 107 => data_o <= "000000000000000000";
        when 108 => data_o <= "000000000000000000";
        when 109 => data_o <= "000000000000000000";
        when 110 => data_o <= "000000000000000000";
        when 111 => data_o <= "000000000000000000";
        when 112 => data_o <= "000000000000000000";
        when 113 => data_o <= "000000000000000000";
        when 114 => data_o <= "000000000000000000";
        when 115 => data_o <= "000000000000000000";
        when 116 => data_o <= "000000000000000000";
        when 117 => data_o <= "000000000000000000";
        when 118 => data_o <= "000000000000000000";
        when 119 => data_o <= "000000000000000000";
        when 120 => data_o <= "000000000000000000";
        when 121 => data_o <= "000000000000000000";
        when 122 => data_o <= "000000000000000000";
        when 123 => data_o <= "000000000000000000";
        when 124 => data_o <= "000000000000000000";
        when 125 => data_o <= "000000000000000000";
        when 126 => data_o <= "000000000000000000";
        when 127 => data_o <= "000000000000000000";
        when 128 => data_o <= "000000000000000000";
        when 129 => data_o <= "000000000000000000";
        when 130 => data_o <= "000000000000000000";
        when 131 => data_o <= "000000000000000000";
        when 132 => data_o <= "000000000000000000";
        when 133 => data_o <= "000000000000000000";
        when 134 => data_o <= "000000000000000000";
        when 135 => data_o <= "000000000000000000";
        when 136 => data_o <= "000000000000000000";
        when 137 => data_o <= "000000000000000000";
        when 138 => data_o <= "000000000000000000";
        when 139 => data_o <= "000000000000000000";
        when 140 => data_o <= "000000000000000000";
        when 141 => data_o <= "000000000000000000";
        when 142 => data_o <= "000000000000000000";
        when 143 => data_o <= "000000000000000000";
        when 144 => data_o <= "000000000000000000";
        when 145 => data_o <= "000000000000000000";
        when 146 => data_o <= "000000000000000000";
        when 147 => data_o <= "000000000000000000";
        when 148 => data_o <= "000000000000000000";
        when 149 => data_o <= "000000000000000000";
        when 150 => data_o <= "000000000000000000";
        when 151 => data_o <= "000000000000000000";
        when 152 => data_o <= "000000000000000000";
        when 153 => data_o <= "000000000000000000";
        when 154 => data_o <= "000000000000000000";
        when 155 => data_o <= "000000000000000000";
        when 156 => data_o <= "000000000000000000";
        when 157 => data_o <= "000000000000000000";
        when 158 => data_o <= "000000000000000000";
        when 159 => data_o <= "000000000000000000";
        when 160 => data_o <= "000000000000000000";
        when 161 => data_o <= "000000000000000000";
        when 162 => data_o <= "000000000000000000";
        when 163 => data_o <= "000000000000000000";
        when 164 => data_o <= "000000000000000000";
        when 165 => data_o <= "000000000000000000";
        when 166 => data_o <= "000000000000000000";
        when 167 => data_o <= "000000000000000000";
        when 168 => data_o <= "000000000000000000";
        when 169 => data_o <= "000000000000000000";
        when 170 => data_o <= "000000000000000000";
        when 171 => data_o <= "000000000000000000";
        when 172 => data_o <= "000000000000000000";
        when 173 => data_o <= "000000000000000000";
        when 174 => data_o <= "000000000000000000";
        when 175 => data_o <= "000000000000000000";
        when 176 => data_o <= "000000000000000000";
        when 177 => data_o <= "000000000000000000";
        when 178 => data_o <= "000000000000000000";
        when 179 => data_o <= "000000000000000000";
        when 180 => data_o <= "000000000000000000";
        when 181 => data_o <= "000000000000000000";
        when 182 => data_o <= "000000000000000000";
        when 183 => data_o <= "000000000000000000";
        when 184 => data_o <= "000000000000000000";
        when 185 => data_o <= "000000000000000000";
        when 186 => data_o <= "000000000000000000";
        when 187 => data_o <= "000000000000000000";
        when 188 => data_o <= "000000000000000000";
        when 189 => data_o <= "000000000000000000";
        when 190 => data_o <= "000000000000000000";
        when 191 => data_o <= "000000000000000000";
        when 192 => data_o <= "000000000000000000";
        when 193 => data_o <= "000000000000000000";
        when 194 => data_o <= "000000000000000000";
        when 195 => data_o <= "000000000000000000";
        when 196 => data_o <= "000000000000000000";
        when 197 => data_o <= "000000000000000000";
        when 198 => data_o <= "000000000000000000";
        when 199 => data_o <= "000000000000000000";
        when 200 => data_o <= "000000000000000000";
        when 201 => data_o <= "000000000000000000";
        when 202 => data_o <= "000000000000000000";
        when 203 => data_o <= "000000000000000000";
        when 204 => data_o <= "000000000000000000";
        when 205 => data_o <= "000000000000000000";
        when 206 => data_o <= "000000000000000000";
        when 207 => data_o <= "000000000000000000";
        when 208 => data_o <= "000000000000000000";
        when 209 => data_o <= "000000000000000000";
        when 210 => data_o <= "000000000000000000";
        when 211 => data_o <= "000000000000000000";
        when 212 => data_o <= "000000000000000000";
        when 213 => data_o <= "000000000000000000";
        when 214 => data_o <= "000000000000000000";
        when 215 => data_o <= "000000000000000000";
        when 216 => data_o <= "000000000000000000";
        when 217 => data_o <= "000000000000000000";
        when 218 => data_o <= "000000000000000000";
        when 219 => data_o <= "000000000000000000";
        when 220 => data_o <= "000000000000000000";
        when 221 => data_o <= "000000000000000000";
        when 222 => data_o <= "000000000000000000";
        when 223 => data_o <= "000000000000000000";
        when 224 => data_o <= "000000000000000000";
        when 225 => data_o <= "000000000000000000";
        when 226 => data_o <= "000000000000000000";
        when 227 => data_o <= "000000000000000000";
        when 228 => data_o <= "000000000000000000";
        when 229 => data_o <= "000000000000000000";
        when 230 => data_o <= "000000000000000000";
        when 231 => data_o <= "000000000000000000";
        when 232 => data_o <= "000000000000000000";
        when 233 => data_o <= "000000000000000000";
        when 234 => data_o <= "000000000000000000";
        when 235 => data_o <= "000000000000000000";
        when 236 => data_o <= "000000000000000000";
        when 237 => data_o <= "000000000000000000";
        when 238 => data_o <= "000000000000000000";
        when 239 => data_o <= "000000000000000000";
        when 240 => data_o <= "000000000000000000";
        when 241 => data_o <= "000000000000000000";
        when 242 => data_o <= "000000000000000000";
        when 243 => data_o <= "000000000000000000";
        when 244 => data_o <= "000000000000000000";
        when 245 => data_o <= "000000000000000000";
        when 246 => data_o <= "000000000000000000";
        when 247 => data_o <= "000000000000000000";
        when 248 => data_o <= "000000000000000000";
        when 249 => data_o <= "000000000000000000";
        when 250 => data_o <= "000000000000000000";
        when 251 => data_o <= "000000000000000000";
        when 252 => data_o <= "000000000000000000";
        when 253 => data_o <= "000000000000000000";
        when 254 => data_o <= "000000000000000000";
        when 255 => data_o <= "000000000000000000";
        when 256 => data_o <= "000000000000000000";
        when 257 => data_o <= "000000000000000000";
        when 258 => data_o <= "000000000000000000";
        when 259 => data_o <= "000000000000000000";
        when 260 => data_o <= "000000000000000000";
        when 261 => data_o <= "000000000000000000";
        when 262 => data_o <= "000000000000000000";
        when 263 => data_o <= "000000000000000000";
        when 264 => data_o <= "000000000000000000";
        when 265 => data_o <= "000000000000000000";
        when 266 => data_o <= "000000000000000000";
        when 267 => data_o <= "000000000000000000";
        when 268 => data_o <= "000000000000000000";
        when 269 => data_o <= "000000000000000000";
        when 270 => data_o <= "000000000000000000";
        when 271 => data_o <= "000000000000000000";
        when 272 => data_o <= "000000000000000000";
        when 273 => data_o <= "000000000000000000";
        when 274 => data_o <= "000000000000000000";
        when 275 => data_o <= "000000000000000000";
        when 276 => data_o <= "000000000000000000";
        when 277 => data_o <= "000000000000000000";
        when 278 => data_o <= "000000000000000000";
        when 279 => data_o <= "000000000000000000";
        when 280 => data_o <= "000000000000000000";
        when 281 => data_o <= "000000000000000000";
        when 282 => data_o <= "000000000000000000";
        when 283 => data_o <= "000000000000000000";
        when 284 => data_o <= "000000000000000000";
        when 285 => data_o <= "000000000000000000";
        when 286 => data_o <= "000000000000000000";
        when 287 => data_o <= "000000000000000000";
        when 288 => data_o <= "000000000000000000";
        when 289 => data_o <= "000000000000000000";
        when 290 => data_o <= "000000000000000000";
        when 291 => data_o <= "000000000000000000";
        when 292 => data_o <= "000000000000000000";
        when 293 => data_o <= "000000000000000000";
        when 294 => data_o <= "000000000000000000";
        when 295 => data_o <= "000000000000000000";
        when 296 => data_o <= "000000000000000000";
        when 297 => data_o <= "000000000000000000";
        when 298 => data_o <= "000000000000000000";
        when 299 => data_o <= "000000000000000000";
        when 300 => data_o <= "000000000000000000";
        when 301 => data_o <= "000000000000000000";
        when 302 => data_o <= "000000000000000000";
        when 303 => data_o <= "000000000000000000";
        when 304 => data_o <= "000000000000000000";
        when 305 => data_o <= "000000000000000000";
        when 306 => data_o <= "000000000000000000";
        when 307 => data_o <= "000000000000000000";
        when 308 => data_o <= "000000000000000000";
        when 309 => data_o <= "000000000000000000";
        when 310 => data_o <= "000000000000000000";
        when 311 => data_o <= "000000000000000000";
        when 312 => data_o <= "000000000000000000";
        when 313 => data_o <= "000000000000000000";
        when 314 => data_o <= "000000000000000000";
        when 315 => data_o <= "000000000000000000";
        when 316 => data_o <= "000000000000000000";
        when 317 => data_o <= "000000000000000000";
        when 318 => data_o <= "000000000000000000";
        when 319 => data_o <= "000000000000000000";
        when 320 => data_o <= "000000000000000000";
        when 321 => data_o <= "000000000000000000";
        when 322 => data_o <= "000000000000000000";
        when 323 => data_o <= "000000000000000000";
        when 324 => data_o <= "000000000000000000";
        when 325 => data_o <= "000000000000000000";
        when 326 => data_o <= "000000000000000000";
        when 327 => data_o <= "000000000000000000";
        when 328 => data_o <= "000000000000000000";
        when 329 => data_o <= "000000000000000000";
        when 330 => data_o <= "000000000000000000";
        when 331 => data_o <= "000000000000000000";
        when 332 => data_o <= "000000000000000000";
        when 333 => data_o <= "000000000000000000";
        when 334 => data_o <= "000000000000000000";
        when 335 => data_o <= "000000000000000000";
        when 336 => data_o <= "000000000000000000";
        when 337 => data_o <= "000000000000000000";
        when 338 => data_o <= "000000000000000000";
        when 339 => data_o <= "000000000000000000";
        when 340 => data_o <= "000000000000000000";
        when 341 => data_o <= "000000000000000000";
        when 342 => data_o <= "000000000000000000";
        when 343 => data_o <= "000000000000000000";
        when 344 => data_o <= "000000000000000000";
        when 345 => data_o <= "000000000000000000";
        when 346 => data_o <= "000000000000000000";
        when 347 => data_o <= "000000000000000000";
        when 348 => data_o <= "000000000000000000";
        when 349 => data_o <= "000000000000000000";
        when 350 => data_o <= "000000000000000000";
        when 351 => data_o <= "000000000000000000";
        when 352 => data_o <= "000000000000000000";
        when 353 => data_o <= "000000000000000000";
        when 354 => data_o <= "000000000000000000";
        when 355 => data_o <= "000000000000000000";
        when 356 => data_o <= "000000000000000000";
        when 357 => data_o <= "000000000000000000";
        when 358 => data_o <= "000000000000000000";
        when 359 => data_o <= "000000000000000000";
        when 360 => data_o <= "000000000000000000";
        when 361 => data_o <= "000000000000000000";
        when 362 => data_o <= "000000000000000000";
        when 363 => data_o <= "000000000000000000";
        when 364 => data_o <= "000000000000000000";
        when 365 => data_o <= "000000000000000000";
        when 366 => data_o <= "000000000000000000";
        when 367 => data_o <= "000000000000000000";
        when 368 => data_o <= "000000000000000000";
        when 369 => data_o <= "000000000000000000";
        when 370 => data_o <= "000000000000000000";
        when 371 => data_o <= "000000000000000000";
        when 372 => data_o <= "000000000000000000";
        when 373 => data_o <= "000000000000000000";
        when 374 => data_o <= "000000000000000000";
        when 375 => data_o <= "000000000000000000";
        when 376 => data_o <= "000000000000000000";
        when 377 => data_o <= "000000000000000000";
        when 378 => data_o <= "000000000000000000";
        when 379 => data_o <= "000000000000000000";
        when 380 => data_o <= "000000000000000000";
        when 381 => data_o <= "000000000000000000";
        when 382 => data_o <= "000000000000000000";
        when 383 => data_o <= "000000000000000000";
        when 384 => data_o <= "000000000000000000";
        when 385 => data_o <= "000000000000000000";
        when 386 => data_o <= "000000000000000000";
        when 387 => data_o <= "000000000000000000";
        when 388 => data_o <= "000000000000000000";
        when 389 => data_o <= "000000000000000000";
        when 390 => data_o <= "000000000000000000";
        when 391 => data_o <= "000000000000000000";
        when 392 => data_o <= "000000000000000000";
        when 393 => data_o <= "000000000000000000";
        when 394 => data_o <= "000000000000000000";
        when 395 => data_o <= "000000000000000000";
        when 396 => data_o <= "000000000000000000";
        when 397 => data_o <= "000000000000000000";
        when 398 => data_o <= "000000000000000000";
        when 399 => data_o <= "000000000000000000";
        when 400 => data_o <= "000000000000000000";
        when 401 => data_o <= "000000000000000000";
        when 402 => data_o <= "000000000000000000";
        when 403 => data_o <= "000000000000000000";
        when 404 => data_o <= "000000000000000000";
        when 405 => data_o <= "000000000000000000";
        when 406 => data_o <= "000000000000000000";
        when 407 => data_o <= "000000000000000000";
        when 408 => data_o <= "000000000000000000";
        when 409 => data_o <= "000000000000000000";
        when 410 => data_o <= "000000000000000000";
        when 411 => data_o <= "000000000000000000";
        when 412 => data_o <= "000000000000000000";
        when 413 => data_o <= "000000000000000000";
        when 414 => data_o <= "000000000000000000";
        when 415 => data_o <= "000000000000000000";
        when 416 => data_o <= "000000000000000000";
        when 417 => data_o <= "000000000000000000";
        when 418 => data_o <= "000000000000000000";
        when 419 => data_o <= "000000000000000000";
        when 420 => data_o <= "000000000000000000";
        when 421 => data_o <= "000000000000000000";
        when 422 => data_o <= "000000000000000000";
        when 423 => data_o <= "000000000000000000";
        when 424 => data_o <= "000000000000000000";
        when 425 => data_o <= "000000000000000000";
        when 426 => data_o <= "000000000000000000";
        when 427 => data_o <= "000000000000000000";
        when 428 => data_o <= "000000000000000000";
        when 429 => data_o <= "000000000000000000";
        when 430 => data_o <= "000000000000000000";
        when 431 => data_o <= "000000000000000000";
        when 432 => data_o <= "000000000000000000";
        when 433 => data_o <= "000000000000000000";
        when 434 => data_o <= "000000000000000000";
        when 435 => data_o <= "000000000000000000";
        when 436 => data_o <= "000000000000000000";
        when 437 => data_o <= "000000000000000000";
        when 438 => data_o <= "000000000000000000";
        when 439 => data_o <= "000000000000000000";
        when 440 => data_o <= "000000000000000000";
        when 441 => data_o <= "000000000000000000";
        when 442 => data_o <= "000000000000000000";
        when 443 => data_o <= "000000000000000000";
        when 444 => data_o <= "000000000000000000";
        when 445 => data_o <= "000000000000000000";
        when 446 => data_o <= "000000000000000000";
        when 447 => data_o <= "000000000000000000";
        when 448 => data_o <= "000000000000000000";
        when 449 => data_o <= "000000000000000000";
        when 450 => data_o <= "000000000000000000";
        when 451 => data_o <= "000000000000000000";
        when 452 => data_o <= "000000000000000000";
        when 453 => data_o <= "000000000000000000";
        when 454 => data_o <= "000000000000000000";
        when 455 => data_o <= "000000000000000000";
        when 456 => data_o <= "000000000000000000";
        when 457 => data_o <= "000000000000000000";
        when 458 => data_o <= "000000000000000000";
        when 459 => data_o <= "000000000000000000";
        when 460 => data_o <= "000000000000000000";
        when 461 => data_o <= "000000000000000000";
        when 462 => data_o <= "000000000000000000";
        when 463 => data_o <= "000000000000000000";
        when 464 => data_o <= "000000000000000000";
        when 465 => data_o <= "000000000000000000";
        when 466 => data_o <= "000000000000000000";
        when 467 => data_o <= "000000000000000000";
        when 468 => data_o <= "000000000000000000";
        when 469 => data_o <= "000000000000000000";
        when 470 => data_o <= "000000000000000000";
        when 471 => data_o <= "000000000000000000";
        when 472 => data_o <= "000000000000000000";
        when 473 => data_o <= "000000000000000000";
        when 474 => data_o <= "000000000000000000";
        when 475 => data_o <= "000000000000000000";
        when 476 => data_o <= "000000000000000000";
        when 477 => data_o <= "000000000000000000";
        when 478 => data_o <= "000000000000000000";
        when 479 => data_o <= "000000000000000000";
        when 480 => data_o <= "000000000000000000";
        when 481 => data_o <= "000000000000000000";
        when 482 => data_o <= "000000000000000000";
        when 483 => data_o <= "000000000000000000";
        when 484 => data_o <= "000000000000000000";
        when 485 => data_o <= "000000000000000000";
        when 486 => data_o <= "000000000000000000";
        when 487 => data_o <= "000000000000000000";
        when 488 => data_o <= "000000000000000000";
        when 489 => data_o <= "000000000000000000";
        when 490 => data_o <= "000000000000000000";
        when 491 => data_o <= "000000000000000000";
        when 492 => data_o <= "000000000000000000";
        when 493 => data_o <= "000000000000000000";
        when 494 => data_o <= "000000000000000000";
        when 495 => data_o <= "000000000000000000";
        when 496 => data_o <= "000000000000000000";
        when 497 => data_o <= "000000000000000000";
        when 498 => data_o <= "000000000000000000";
        when 499 => data_o <= "000000000000000000";
        when 500 => data_o <= "000000000000000000";
        when 501 => data_o <= "000000000000000000";
        when 502 => data_o <= "000000000000000000";
        when 503 => data_o <= "000000000000000000";
        when 504 => data_o <= "000000000000000000";
        when 505 => data_o <= "000000000000000000";
        when 506 => data_o <= "000000000000000000";
        when 507 => data_o <= "000000000000000000";
        when 508 => data_o <= "000000000000000000";
        when 509 => data_o <= "000000000000000000";
        when 510 => data_o <= "000000000000000000";
        when 511 => data_o <= "000000000000000000";
        when 512 => data_o <= "000000000000000000";
        when 513 => data_o <= "000000000000000000";
        when 514 => data_o <= "000000000000000000";
        when 515 => data_o <= "000000000000000000";
        when 516 => data_o <= "000000000000000000";
        when 517 => data_o <= "000000000000000000";
        when 518 => data_o <= "000000000000000000";
        when 519 => data_o <= "000000000000000000";
        when 520 => data_o <= "000000000000000000";
        when 521 => data_o <= "000000000000000000";
        when 522 => data_o <= "000000000000000000";
        when 523 => data_o <= "000000000000000000";
        when 524 => data_o <= "000000000000000000";
        when 525 => data_o <= "000000000000000000";
        when 526 => data_o <= "000000000000000000";
        when 527 => data_o <= "000000000000000000";
        when 528 => data_o <= "000000000000000000";
        when 529 => data_o <= "000000000000000000";
        when 530 => data_o <= "000000000000000000";
        when 531 => data_o <= "000000000000000000";
        when 532 => data_o <= "000000000000000000";
        when 533 => data_o <= "000000000000000000";
        when 534 => data_o <= "000000000000000000";
        when 535 => data_o <= "000000000000000000";
        when 536 => data_o <= "000000000000000000";
        when 537 => data_o <= "000000000000000000";
        when 538 => data_o <= "000000000000000000";
        when 539 => data_o <= "000000000000000000";
        when 540 => data_o <= "000000000000000000";
        when 541 => data_o <= "000000000000000000";
        when 542 => data_o <= "000000000000000000";
        when 543 => data_o <= "000000000000000000";
        when 544 => data_o <= "000000000000000000";
        when 545 => data_o <= "000000000000000000";
        when 546 => data_o <= "000000000000000000";
        when 547 => data_o <= "000000000000000000";
        when 548 => data_o <= "000000000000000000";
        when 549 => data_o <= "000000000000000000";
        when 550 => data_o <= "000000000000000000";
        when 551 => data_o <= "000000000000000000";
        when 552 => data_o <= "000000000000000000";
        when 553 => data_o <= "000000000000000000";
        when 554 => data_o <= "000000000000000000";
        when 555 => data_o <= "000000000000000000";
        when 556 => data_o <= "000000000000000000";
        when 557 => data_o <= "000000000000000000";
        when 558 => data_o <= "000000000000000000";
        when 559 => data_o <= "000000000000000000";
        when 560 => data_o <= "000000000000000000";
        when 561 => data_o <= "000000000000000000";
        when 562 => data_o <= "000000000000000000";
        when 563 => data_o <= "000000000000000000";
        when 564 => data_o <= "000000000000000000";
        when 565 => data_o <= "000000000000000000";
        when 566 => data_o <= "000000000000000000";
        when 567 => data_o <= "000000000000000000";
        when 568 => data_o <= "000000000000000000";
        when 569 => data_o <= "000000000000000000";
        when 570 => data_o <= "000000000000000000";
        when 571 => data_o <= "000000000000000000";
        when 572 => data_o <= "000000000000000000";
        when 573 => data_o <= "000000000000000000";
        when 574 => data_o <= "000000000000000000";
        when 575 => data_o <= "000000000000000000";
        when 576 => data_o <= "000000000000000000";
        when 577 => data_o <= "000000000000000000";
        when 578 => data_o <= "000000000000000000";
        when 579 => data_o <= "000000000000000000";
        when 580 => data_o <= "000000000000000000";
        when 581 => data_o <= "000000000000000000";
        when 582 => data_o <= "000000000000000000";
        when 583 => data_o <= "000000000000000000";
        when 584 => data_o <= "000000000000000000";
        when 585 => data_o <= "000000000000000000";
        when 586 => data_o <= "000000000000000000";
        when 587 => data_o <= "000000000000000000";
        when 588 => data_o <= "000000000000000000";
        when 589 => data_o <= "000000000000000000";
        when 590 => data_o <= "000000000000000000";
        when 591 => data_o <= "000000000000000000";
        when 592 => data_o <= "000000000000000000";
        when 593 => data_o <= "000000000000000000";
        when 594 => data_o <= "000000000000000000";
        when 595 => data_o <= "000000000000000000";
        when 596 => data_o <= "000000000000000000";
        when 597 => data_o <= "000000000000000000";
        when 598 => data_o <= "000000000000000000";
        when 599 => data_o <= "000000000000000000";
        when 600 => data_o <= "000000000000000000";
        when 601 => data_o <= "000000000000000000";
        when 602 => data_o <= "000000000000000000";
        when 603 => data_o <= "000000000000000000";
        when 604 => data_o <= "000000000000000000";
        when 605 => data_o <= "000000000000000000";
        when 606 => data_o <= "000000000000000000";
        when 607 => data_o <= "000000000000000000";
        when 608 => data_o <= "000000000000000000";
        when 609 => data_o <= "000000000000000000";
        when 610 => data_o <= "000000000000000000";
        when 611 => data_o <= "000000000000000000";
        when 612 => data_o <= "000000000000000000";
        when 613 => data_o <= "000000000000000000";
        when 614 => data_o <= "000000000000000000";
        when 615 => data_o <= "000000000000000000";
        when 616 => data_o <= "000000000000000000";
        when 617 => data_o <= "000000000000000000";
        when 618 => data_o <= "000000000000000000";
        when 619 => data_o <= "000000000000000000";
        when 620 => data_o <= "000000000000000000";
        when 621 => data_o <= "000000000000000000";
        when 622 => data_o <= "000000000000000000";
        when 623 => data_o <= "000000000000000000";
        when 624 => data_o <= "000000000000000000";
        when 625 => data_o <= "000000000000000000";
        when 626 => data_o <= "000000000000000000";
        when 627 => data_o <= "000000000000000000";
        when 628 => data_o <= "000000000000000000";
        when 629 => data_o <= "000000000000000000";
        when 630 => data_o <= "000000000000000000";
        when 631 => data_o <= "000000000000000000";
        when 632 => data_o <= "000000000000000000";
        when 633 => data_o <= "000000000000000000";
        when 634 => data_o <= "000000000000000000";
        when 635 => data_o <= "000000000000000000";
        when 636 => data_o <= "000000000000000000";
        when 637 => data_o <= "000000000000000000";
        when 638 => data_o <= "000000000000000000";
        when 639 => data_o <= "000000000000000000";
        when 640 => data_o <= "000000000000000000";
        when 641 => data_o <= "000000000000000000";
        when 642 => data_o <= "000000000000000000";
        when 643 => data_o <= "000000000000000000";
        when 644 => data_o <= "000000000000000000";
        when 645 => data_o <= "000000000000000000";
        when 646 => data_o <= "000000000000000000";
        when 647 => data_o <= "000000000000000000";
        when 648 => data_o <= "000000000000000000";
        when 649 => data_o <= "000000000000000000";
        when 650 => data_o <= "000000000000000000";
        when 651 => data_o <= "000000000000000000";
        when 652 => data_o <= "000000000000000000";
        when 653 => data_o <= "000000000000000000";
        when 654 => data_o <= "000000000000000000";
        when 655 => data_o <= "000000000000000000";
        when 656 => data_o <= "000000000000000000";
        when 657 => data_o <= "000000000000000000";
        when 658 => data_o <= "000000000000000000";
        when 659 => data_o <= "000000000000000000";
        when 660 => data_o <= "000000000000000000";
        when 661 => data_o <= "000000000000000000";
        when 662 => data_o <= "000000000000000000";
        when 663 => data_o <= "000000000000000000";
        when 664 => data_o <= "000000000000000000";
        when 665 => data_o <= "000000000000000000";
        when 666 => data_o <= "000000000000000000";
        when 667 => data_o <= "000000000000000000";
        when 668 => data_o <= "000000000000000000";
        when 669 => data_o <= "000000000000000000";
        when 670 => data_o <= "000000000000000000";
        when 671 => data_o <= "000000000000000000";
        when 672 => data_o <= "000000000000000000";
        when 673 => data_o <= "000000000000000000";
        when 674 => data_o <= "000000000000000000";
        when 675 => data_o <= "000000000000000000";
        when 676 => data_o <= "000000000000000000";
        when 677 => data_o <= "000000000000000000";
        when 678 => data_o <= "000000000000000000";
        when 679 => data_o <= "000000000000000000";
        when 680 => data_o <= "000000000000000000";
        when 681 => data_o <= "000000000000000000";
        when 682 => data_o <= "000000000000000000";
        when 683 => data_o <= "000000000000000000";
        when 684 => data_o <= "000000000000000000";
        when 685 => data_o <= "000000000000000000";
        when 686 => data_o <= "000000000000000000";
        when 687 => data_o <= "000000000000000000";
        when 688 => data_o <= "000000000000000000";
        when 689 => data_o <= "000000000000000000";
        when 690 => data_o <= "000000000000000000";
        when 691 => data_o <= "000000000000000000";
        when 692 => data_o <= "000000000000000000";
        when 693 => data_o <= "000000000000000000";
        when 694 => data_o <= "000000000000000000";
        when 695 => data_o <= "000000000000000000";
        when 696 => data_o <= "000000000000000000";
        when 697 => data_o <= "000000000000000000";
        when 698 => data_o <= "000000000000000000";
        when 699 => data_o <= "000000000000000000";
        when 700 => data_o <= "000000000000000000";
        when 701 => data_o <= "000000000000000000";
        when 702 => data_o <= "000000000000000000";
        when 703 => data_o <= "000000000000000000";
        when 704 => data_o <= "000000000000000000";
        when 705 => data_o <= "000000000000000000";
        when 706 => data_o <= "000000000000000000";
        when 707 => data_o <= "000000000000000000";
        when 708 => data_o <= "000000000000000000";
        when 709 => data_o <= "000000000000000000";
        when 710 => data_o <= "000000000000000000";
        when 711 => data_o <= "000000000000000000";
        when 712 => data_o <= "000000000000000000";
        when 713 => data_o <= "000000000000000000";
        when 714 => data_o <= "000000000000000000";
        when 715 => data_o <= "000000000000000000";
        when 716 => data_o <= "000000000000000000";
        when 717 => data_o <= "000000000000000000";
        when 718 => data_o <= "000000000000000000";
        when 719 => data_o <= "000000000000000000";
        when 720 => data_o <= "000000000000000000";
        when 721 => data_o <= "000000000000000000";
        when 722 => data_o <= "000000000000000000";
        when 723 => data_o <= "000000000000000000";
        when 724 => data_o <= "000000000000000000";
        when 725 => data_o <= "000000000000000000";
        when 726 => data_o <= "000000000000000000";
        when 727 => data_o <= "000000000000000000";
        when 728 => data_o <= "000000000000000000";
        when 729 => data_o <= "000000000000000000";
        when 730 => data_o <= "000000000000000000";
        when 731 => data_o <= "000000000000000000";
        when 732 => data_o <= "000000000000000000";
        when 733 => data_o <= "000000000000000000";
        when 734 => data_o <= "000000000000000000";
        when 735 => data_o <= "000000000000000000";
        when 736 => data_o <= "000000000000000000";
        when 737 => data_o <= "000000000000000000";
        when 738 => data_o <= "000000000000000000";
        when 739 => data_o <= "000000000000000000";
        when 740 => data_o <= "000000000000000000";
        when 741 => data_o <= "000000000000000000";
        when 742 => data_o <= "000000000000000000";
        when 743 => data_o <= "000000000000000000";
        when 744 => data_o <= "000000000000000000";
        when 745 => data_o <= "000000000000000000";
        when 746 => data_o <= "000000000000000000";
        when 747 => data_o <= "000000000000000000";
        when 748 => data_o <= "000000000000000000";
        when 749 => data_o <= "000000000000000000";
        when 750 => data_o <= "000000000000000000";
        when 751 => data_o <= "000000000000000000";
        when 752 => data_o <= "000000000000000000";
        when 753 => data_o <= "000000000000000000";
        when 754 => data_o <= "000000000000000000";
        when 755 => data_o <= "000000000000000000";
        when 756 => data_o <= "000000000000000000";
        when 757 => data_o <= "000000000000000000";
        when 758 => data_o <= "000000000000000000";
        when 759 => data_o <= "000000000000000000";
        when 760 => data_o <= "000000000000000000";
        when 761 => data_o <= "000000000000000000";
        when 762 => data_o <= "000000000000000000";
        when 763 => data_o <= "000000000000000000";
        when 764 => data_o <= "000000000000000000";
        when 765 => data_o <= "000000000000000000";
        when 766 => data_o <= "000000000000000000";
        when 767 => data_o <= "000000000000000000";
        when 768 => data_o <= "000000000000000000";
        when 769 => data_o <= "000000000000000000";
        when 770 => data_o <= "000000000000000000";
        when 771 => data_o <= "000000000000000000";
        when 772 => data_o <= "000000000000000000";
        when 773 => data_o <= "000000000000000000";
        when 774 => data_o <= "000000000000000000";
        when 775 => data_o <= "000000000000000000";
        when 776 => data_o <= "000000000000000000";
        when 777 => data_o <= "000000000000000000";
        when 778 => data_o <= "000000000000000000";
        when 779 => data_o <= "000000000000000000";
        when 780 => data_o <= "000000000000000000";
        when 781 => data_o <= "000000000000000000";
        when 782 => data_o <= "000000000000000000";
        when 783 => data_o <= "000000000000000000";
        when 784 => data_o <= "000000000000000000";
        when 785 => data_o <= "000000000000000000";
        when 786 => data_o <= "000000000000000000";
        when 787 => data_o <= "000000000000000000";
        when 788 => data_o <= "000000000000000000";
        when 789 => data_o <= "000000000000000000";
        when 790 => data_o <= "000000000000000000";
        when 791 => data_o <= "000000000000000000";
        when 792 => data_o <= "000000000000000000";
        when 793 => data_o <= "000000000000000000";
        when 794 => data_o <= "000000000000000000";
        when 795 => data_o <= "000000000000000000";
        when 796 => data_o <= "000000000000000000";
        when 797 => data_o <= "000000000000000000";
        when 798 => data_o <= "000000000000000000";
        when 799 => data_o <= "000000000000000000";
        when 800 => data_o <= "000000000000000000";
        when 801 => data_o <= "000000000000000000";
        when 802 => data_o <= "000000000000000000";
        when 803 => data_o <= "000000000000000000";
        when 804 => data_o <= "000000000000000000";
        when 805 => data_o <= "000000000000000000";
        when 806 => data_o <= "000000000000000000";
        when 807 => data_o <= "000000000000000000";
        when 808 => data_o <= "000000000000000000";
        when 809 => data_o <= "000000000000000000";
        when 810 => data_o <= "000000000000000000";
        when 811 => data_o <= "000000000000000000";
        when 812 => data_o <= "000000000000000000";
        when 813 => data_o <= "000000000000000000";
        when 814 => data_o <= "000000000000000000";
        when 815 => data_o <= "000000000000000000";
        when 816 => data_o <= "000000000000000000";
        when 817 => data_o <= "000000000000000000";
        when 818 => data_o <= "000000000000000000";
        when 819 => data_o <= "000000000000000000";
        when 820 => data_o <= "000000000000000000";
        when 821 => data_o <= "000000000000000000";
        when 822 => data_o <= "000000000000000000";
        when 823 => data_o <= "000000000000000000";
        when 824 => data_o <= "000000000000000000";
        when 825 => data_o <= "000000000000000000";
        when 826 => data_o <= "000000000000000000";
        when 827 => data_o <= "000000000000000000";
        when 828 => data_o <= "000000000000000000";
        when 829 => data_o <= "000000000000000000";
        when 830 => data_o <= "000000000000000000";
        when 831 => data_o <= "000000000000000000";
        when 832 => data_o <= "000000000000000000";
        when 833 => data_o <= "000000000000000000";
        when 834 => data_o <= "000000000000000000";
        when 835 => data_o <= "000000000000000000";
        when 836 => data_o <= "000000000000000000";
        when 837 => data_o <= "000000000000000000";
        when 838 => data_o <= "000000000000000000";
        when 839 => data_o <= "000000000000000000";
        when 840 => data_o <= "000000000000000000";
        when 841 => data_o <= "000000000000000000";
        when 842 => data_o <= "000000000000000000";
        when 843 => data_o <= "000000000000000000";
        when 844 => data_o <= "000000000000000000";
        when 845 => data_o <= "000000000000000000";
        when 846 => data_o <= "000000000000000000";
        when 847 => data_o <= "000000000000000000";
        when 848 => data_o <= "000000000000000000";
        when 849 => data_o <= "000000000000000000";
        when 850 => data_o <= "000000000000000000";
        when 851 => data_o <= "000000000000000000";
        when 852 => data_o <= "000000000000000000";
        when 853 => data_o <= "000000000000000000";
        when 854 => data_o <= "000000000000000000";
        when 855 => data_o <= "000000000000000000";
        when 856 => data_o <= "000000000000000000";
        when 857 => data_o <= "000000000000000000";
        when 858 => data_o <= "000000000000000000";
        when 859 => data_o <= "000000000000000000";
        when 860 => data_o <= "000000000000000000";
        when 861 => data_o <= "000000000000000000";
        when 862 => data_o <= "000000000000000000";
        when 863 => data_o <= "000000000000000000";
        when 864 => data_o <= "000000000000000000";
        when 865 => data_o <= "000000000000000000";
        when 866 => data_o <= "000000000000000000";
        when 867 => data_o <= "000000000000000000";
        when 868 => data_o <= "000000000000000000";
        when 869 => data_o <= "000000000000000000";
        when 870 => data_o <= "000000000000000000";
        when 871 => data_o <= "000000000000000000";
        when 872 => data_o <= "000000000000000000";
        when 873 => data_o <= "000000000000000000";
        when 874 => data_o <= "000000000000000000";
        when 875 => data_o <= "000000000000000000";
        when 876 => data_o <= "000000000000000000";
        when 877 => data_o <= "000000000000000000";
        when 878 => data_o <= "000000000000000000";
        when 879 => data_o <= "000000000000000000";
        when 880 => data_o <= "000000000000000000";
        when 881 => data_o <= "000000000000000000";
        when 882 => data_o <= "000000000000000000";
        when 883 => data_o <= "000000000000000000";
        when 884 => data_o <= "000000000000000000";
        when 885 => data_o <= "000000000000000000";
        when 886 => data_o <= "000000000000000000";
        when 887 => data_o <= "000000000000000000";
        when 888 => data_o <= "000000000000000000";
        when 889 => data_o <= "000000000000000000";
        when 890 => data_o <= "000000000000000000";
        when 891 => data_o <= "000000000000000000";
        when 892 => data_o <= "000000000000000000";
        when 893 => data_o <= "000000000000000000";
        when 894 => data_o <= "000000000000000000";
        when 895 => data_o <= "000000000000000000";
        when 896 => data_o <= "000000000000000000";
        when 897 => data_o <= "000000000000000000";
        when 898 => data_o <= "000000000000000000";
        when 899 => data_o <= "000000000000000000";
        when 900 => data_o <= "000000000000000000";
        when 901 => data_o <= "000000000000000000";
        when 902 => data_o <= "000000000000000000";
        when 903 => data_o <= "000000000000000000";
        when 904 => data_o <= "000000000000000000";
        when 905 => data_o <= "000000000000000000";
        when 906 => data_o <= "000000000000000000";
        when 907 => data_o <= "000000000000000000";
        when 908 => data_o <= "000000000000000000";
        when 909 => data_o <= "000000000000000000";
        when 910 => data_o <= "000000000000000000";
        when 911 => data_o <= "000000000000000000";
        when 912 => data_o <= "000000000000000000";
        when 913 => data_o <= "000000000000000000";
        when 914 => data_o <= "000000000000000000";
        when 915 => data_o <= "000000000000000000";
        when 916 => data_o <= "000000000000000000";
        when 917 => data_o <= "000000000000000000";
        when 918 => data_o <= "000000000000000000";
        when 919 => data_o <= "000000000000000000";
        when 920 => data_o <= "000000000000000000";
        when 921 => data_o <= "000000000000000000";
        when 922 => data_o <= "000000000000000000";
        when 923 => data_o <= "000000000000000000";
        when 924 => data_o <= "000000000000000000";
        when 925 => data_o <= "000000000000000000";
        when 926 => data_o <= "000000000000000000";
        when 927 => data_o <= "000000000000000000";
        when 928 => data_o <= "000000000000000000";
        when 929 => data_o <= "000000000000000000";
        when 930 => data_o <= "000000000000000000";
        when 931 => data_o <= "000000000000000000";
        when 932 => data_o <= "000000000000000000";
        when 933 => data_o <= "000000000000000000";
        when 934 => data_o <= "000000000000000000";
        when 935 => data_o <= "000000000000000000";
        when 936 => data_o <= "000000000000000000";
        when 937 => data_o <= "000000000000000000";
        when 938 => data_o <= "000000000000000000";
        when 939 => data_o <= "000000000000000000";
        when 940 => data_o <= "000000000000000000";
        when 941 => data_o <= "000000000000000000";
        when 942 => data_o <= "000000000000000000";
        when 943 => data_o <= "000000000000000000";
        when 944 => data_o <= "000000000000000000";
        when 945 => data_o <= "000000000000000000";
        when 946 => data_o <= "000000000000000000";
        when 947 => data_o <= "000000000000000000";
        when 948 => data_o <= "000000000000000000";
        when 949 => data_o <= "000000000000000000";
        when 950 => data_o <= "000000000000000000";
        when 951 => data_o <= "000000000000000000";
        when 952 => data_o <= "000000000000000000";
        when 953 => data_o <= "000000000000000000";
        when 954 => data_o <= "000000000000000000";
        when 955 => data_o <= "000000000000000000";
        when 956 => data_o <= "000000000000000000";
        when 957 => data_o <= "000000000000000000";
        when 958 => data_o <= "000000000000000000";
        when 959 => data_o <= "000000000000000000";
        when 960 => data_o <= "000000000000000000";
        when 961 => data_o <= "000000000000000000";
        when 962 => data_o <= "000000000000000000";
        when 963 => data_o <= "000000000000000000";
        when 964 => data_o <= "000000000000000000";
        when 965 => data_o <= "000000000000000000";
        when 966 => data_o <= "000000000000000000";
        when 967 => data_o <= "000000000000000000";
        when 968 => data_o <= "000000000000000000";
        when 969 => data_o <= "000000000000000000";
        when 970 => data_o <= "000000000000000000";
        when 971 => data_o <= "000000000000000000";
        when 972 => data_o <= "000000000000000000";
        when 973 => data_o <= "000000000000000000";
        when 974 => data_o <= "000000000000000000";
        when 975 => data_o <= "000000000000000000";
        when 976 => data_o <= "000000000000000000";
        when 977 => data_o <= "000000000000000000";
        when 978 => data_o <= "000000000000000000";
        when 979 => data_o <= "000000000000000000";
        when 980 => data_o <= "000000000000000000";
        when 981 => data_o <= "000000000000000000";
        when 982 => data_o <= "000000000000000000";
        when 983 => data_o <= "000000000000000000";
        when 984 => data_o <= "000000000000000000";
        when 985 => data_o <= "000000000000000000";
        when 986 => data_o <= "000000000000000000";
        when 987 => data_o <= "000000000000000000";
        when 988 => data_o <= "000000000000000000";
        when 989 => data_o <= "000000000000000000";
        when 990 => data_o <= "000000000000000000";
        when 991 => data_o <= "000000000000000000";
        when 992 => data_o <= "000000000000000000";
        when 993 => data_o <= "000000000000000000";
        when 994 => data_o <= "000000000000000000";
        when 995 => data_o <= "000000000000000000";
        when 996 => data_o <= "000000000000000000";
        when 997 => data_o <= "000000000000000000";
        when 998 => data_o <= "000000000000000000";
        when 999 => data_o <= "000000000000000000";
        when 1000 => data_o <= "000000000000000000";
        when 1001 => data_o <= "000000000000000000";
        when 1002 => data_o <= "000000000000000000";
        when 1003 => data_o <= "000000000000000000";
        when 1004 => data_o <= "000000000000000000";
        when 1005 => data_o <= "000000000000000000";
        when 1006 => data_o <= "000000000000000000";
        when 1007 => data_o <= "000000000000000000";
        when 1008 => data_o <= "000000000000000000";
        when 1009 => data_o <= "000000000000000000";
        when 1010 => data_o <= "000000000000000000";
        when 1011 => data_o <= "000000000000000000";
        when 1012 => data_o <= "000000000000000000";
        when 1013 => data_o <= "000000000000000000";
        when 1014 => data_o <= "000000000000000000";
        when 1015 => data_o <= "000000000000000000";
        when 1016 => data_o <= "000000000000000000";
        when 1017 => data_o <= "000000000000000000";
        when 1018 => data_o <= "000000000000000000";
        when 1019 => data_o <= "000000000000000000";
        when 1020 => data_o <= "000000000000000000";
        when 1021 => data_o <= "000000000000000000";
        when 1022 => data_o <= "000000000000000000";
        when 1023 => data_o <= "111000000000000001";
        when others => data_o <= (OTHERS => '0');
      end case;
    end if;
  end process;
end behavioral;
