library IEEE ;
use IEEE.STD_LOGIC_1164.all ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;


entity OpenBlaze8_ROM is   
generic (   ADDRSIZE : natural:=10;      --a modifier 
            INSTSIZE : natural:=18;      --si on change de cible spartan
            JADDRSIZE : natural:=11;     --trois cibles fpga virtex  s2  S3
            JDATASIZE : natural:=9);     -- ou coolruner
    port ( 
        clk_i : in std_logic ;
--      reset : out std_logic ;
        addr_i : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        data_o : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity OpenBlaze8_ROM ;

architecture rtl of OpenBlaze8_ROM is


    component jtag_shifter is
        port ( 
			clk : in std_logic ;
			user1 : out std_logic ;
            write : out std_logic ;
            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
        ) ;
    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18 :  if addrsize /= 0 generate
	    attribute INIT_00 of bram : label is "0066C00A0065C00A0065C00A0062C00A0064C00A0061C00A0065C00A00640E41" ;
	    attribute INIT_01 of bram : label is "002400240024002400240024002440110019EEFFCE09C008C004A0014000C00A" ;
	    attribute INIT_02 of bram : label is "20024010C0100011C0100000C01400648F01F0F0A0000034A000002400240024" ;
	    attribute INIT_03 of bram : label is "404102F7404301774045002A8F01F2F08F01F1F08F01F0F0A00070F0CF01502E" ;
	    attribute INIT_04 of bram : label is "000000000000A00070F0CF0171F0CF0172F0CF01543CC001543EC1015440C201" ;
	    attribute INIT_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_07 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_08 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_09 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_10 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_11 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_12 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_13 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_14 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_15 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_16 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_17 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_18 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_19 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_35 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "8001000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_00 of bram : label is "00000000000000000000000002111DDDCCC6668748886BBFFFFFCA8222222220" ;
	    attribute INITP_01 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_02 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "C000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"0066C00A0065C00A0065C00A0062C00A0064C00A0061C00A0065C00A00640E41",
	            INIT_01 => X"002400240024002400240024002440110019EEFFCE09C008C004A0014000C00A",
	            INIT_02 => X"20024010C0100011C0100000C01400648F01F0F0A0000034A000002400240024",
	            INIT_03 => X"404102F7404301774045002A8F01F2F08F01F1F08F01F0F0A00070F0CF01502E",
	            INIT_04 => X"000000000000A00070F0CF0171F0CF0172F0CF01543CC001543EC1015440C201",
	            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"8001000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"00000000000000000000000002111DDDCCC6668748886BBFFFFFCA8222222220",
	            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )

	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk_i,
	            ADDRB => addr_i,
	            DOB => data_o( 18 - 3 downto 0 ),
	            DOPB => data_o( 18 - 1 downto 18 - 2 ),
	            DIA => jdata( 9 - 2 downto 0 ),
	            DIPA => jdata( 9 - 1 downto 9 - 1 ),
	            ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk_i,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture rtl ;
