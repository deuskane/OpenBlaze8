library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OpenBlaze8_ROM is
  port (
    clk_i    : in std_logic;
    addr_i   : in std_logic_vector(9 downto 0);
    data_o   : out std_logic_vector(17 downto 0)
  );
end OpenBlaze8_ROM ;

architecture rtl of OpenBlaze8_ROM is
  type rom_t is array (0 to 1024-1) of std_logic_vector(18-1 downto 0);
  signal rom : rom_t :=
   (
    0 => "000000111000000000"
   ,1 => "000000000001100100"
   ,2 => "101100000000001010"
   ,3 => "000000000001100101"
   ,4 => "101100000000001010"
   ,5 => "000000000001100001"
   ,6 => "101100000000001010"
   ,7 => "000000000001100100"
   ,8 => "101100000000001010"
   ,9 => "000000000001100010"
   ,10 => "101100000000001010"
   ,11 => "000000000001100101"
   ,12 => "101100000000001010"
   ,13 => "000000000001100101"
   ,14 => "101100000000001010"
   ,15 => "000000000001100110"
   ,16 => "101100000000001010"
   ,17 => "000100000000000000"
   ,18 => "001010000000000001"
   ,19 => "101100000000000100"
   ,20 => "101100000000001000"
   ,21 => "101100111000001001"
   ,22 => "011000111000000001"
   ,23 => "110000000000100100"
   ,24 => "110100000000010001"
   ,25 => "110000000000100100"
   ,26 => "110000000000100100"
   ,27 => "110000000000100100"
   ,28 => "110000000000100100"
   ,29 => "110000000000100100"
   ,30 => "110000000000100100"
   ,31 => "110000000000100100"
   ,32 => "110000000000100100"
   ,33 => "110000000000100100"
   ,34 => "110000000000100100"
   ,35 => "101010000000000000"
   ,36 => "101111000011110000"
   ,37 => "011000111100000001"
   ,38 => "101111000111110000"
   ,39 => "011000111100000001"
   ,40 => "101111001011110000"
   ,41 => "011000111100000001"
   ,42 => "000000000000101010"
   ,43 => "110100000000110101"
   ,44 => "000000000101110111"
   ,45 => "110100000000110011"
   ,46 => "000000001011110111"
   ,47 => "110100000000110001"
   ,48 => "011100001000000001"
   ,49 => "110101010000110000"
   ,50 => "011100000100000001"
   ,51 => "110101010000101110"
   ,52 => "011100000000000001"
   ,53 => "110101010000101100"
   ,54 => "011100111100000001"
   ,55 => "000111001011110000"
   ,56 => "011100111100000001"
   ,57 => "000111000111110000"
   ,58 => "011100111100000001"
   ,59 => "000111000011110000"
   ,60 => "101010000000000000"
   ,61 => "000000000000000000"
   ,62 => "000000000000000000"
   ,63 => "000000000000000000"
   ,64 => "000000000000000000"
   ,65 => "000000000000000000"
   ,66 => "000000000000000000"
   ,67 => "000000000000000000"
   ,68 => "000000000000000000"
   ,69 => "000000000000000000"
   ,70 => "000000000000000000"
   ,71 => "000000000000000000"
   ,72 => "000000000000000000"
   ,73 => "000000000000000000"
   ,74 => "000000000000000000"
   ,75 => "000000000000000000"
   ,76 => "000000000000000000"
   ,77 => "000000000000000000"
   ,78 => "000000000000000000"
   ,79 => "000000000000000000"
   ,80 => "000000000000000000"
   ,81 => "000000000000000000"
   ,82 => "000000000000000000"
   ,83 => "000000000000000000"
   ,84 => "000000000000000000"
   ,85 => "000000000000000000"
   ,86 => "000000000000000000"
   ,87 => "000000000000000000"
   ,88 => "000000000000000000"
   ,89 => "000000000000000000"
   ,90 => "000000000000000000"
   ,91 => "000000000000000000"
   ,92 => "000000000000000000"
   ,93 => "000000000000000000"
   ,94 => "000000000000000000"
   ,95 => "000000000000000000"
   ,96 => "000000000000000000"
   ,97 => "000000000000000000"
   ,98 => "000000000000000000"
   ,99 => "000000000000000000"
   ,100 => "000000000000000000"
   ,101 => "000000000000000000"
   ,102 => "000000000000000000"
   ,103 => "000000000000000000"
   ,104 => "000000000000000000"
   ,105 => "000000000000000000"
   ,106 => "000000000000000000"
   ,107 => "000000000000000000"
   ,108 => "000000000000000000"
   ,109 => "000000000000000000"
   ,110 => "000000000000000000"
   ,111 => "000000000000000000"
   ,112 => "000000000000000000"
   ,113 => "000000000000000000"
   ,114 => "000000000000000000"
   ,115 => "000000000000000000"
   ,116 => "000000000000000000"
   ,117 => "000000000000000000"
   ,118 => "000000000000000000"
   ,119 => "000000000000000000"
   ,120 => "000000000000000000"
   ,121 => "000000000000000000"
   ,122 => "000000000000000000"
   ,123 => "000000000000000000"
   ,124 => "000000000000000000"
   ,125 => "000000000000000000"
   ,126 => "000000000000000000"
   ,127 => "000000000000000000"
   ,128 => "000000000000000000"
   ,129 => "000000000000000000"
   ,130 => "000000000000000000"
   ,131 => "000000000000000000"
   ,132 => "000000000000000000"
   ,133 => "000000000000000000"
   ,134 => "000000000000000000"
   ,135 => "000000000000000000"
   ,136 => "000000000000000000"
   ,137 => "000000000000000000"
   ,138 => "000000000000000000"
   ,139 => "000000000000000000"
   ,140 => "000000000000000000"
   ,141 => "000000000000000000"
   ,142 => "000000000000000000"
   ,143 => "000000000000000000"
   ,144 => "000000000000000000"
   ,145 => "000000000000000000"
   ,146 => "000000000000000000"
   ,147 => "000000000000000000"
   ,148 => "000000000000000000"
   ,149 => "000000000000000000"
   ,150 => "000000000000000000"
   ,151 => "000000000000000000"
   ,152 => "000000000000000000"
   ,153 => "000000000000000000"
   ,154 => "000000000000000000"
   ,155 => "000000000000000000"
   ,156 => "000000000000000000"
   ,157 => "000000000000000000"
   ,158 => "000000000000000000"
   ,159 => "000000000000000000"
   ,160 => "000000000000000000"
   ,161 => "000000000000000000"
   ,162 => "000000000000000000"
   ,163 => "000000000000000000"
   ,164 => "000000000000000000"
   ,165 => "000000000000000000"
   ,166 => "000000000000000000"
   ,167 => "000000000000000000"
   ,168 => "000000000000000000"
   ,169 => "000000000000000000"
   ,170 => "000000000000000000"
   ,171 => "000000000000000000"
   ,172 => "000000000000000000"
   ,173 => "000000000000000000"
   ,174 => "000000000000000000"
   ,175 => "000000000000000000"
   ,176 => "000000000000000000"
   ,177 => "000000000000000000"
   ,178 => "000000000000000000"
   ,179 => "000000000000000000"
   ,180 => "000000000000000000"
   ,181 => "000000000000000000"
   ,182 => "000000000000000000"
   ,183 => "000000000000000000"
   ,184 => "000000000000000000"
   ,185 => "000000000000000000"
   ,186 => "000000000000000000"
   ,187 => "000000000000000000"
   ,188 => "000000000000000000"
   ,189 => "000000000000000000"
   ,190 => "000000000000000000"
   ,191 => "000000000000000000"
   ,192 => "000000000000000000"
   ,193 => "000000000000000000"
   ,194 => "000000000000000000"
   ,195 => "000000000000000000"
   ,196 => "000000000000000000"
   ,197 => "000000000000000000"
   ,198 => "000000000000000000"
   ,199 => "000000000000000000"
   ,200 => "000000000000000000"
   ,201 => "000000000000000000"
   ,202 => "000000000000000000"
   ,203 => "000000000000000000"
   ,204 => "000000000000000000"
   ,205 => "000000000000000000"
   ,206 => "000000000000000000"
   ,207 => "000000000000000000"
   ,208 => "000000000000000000"
   ,209 => "000000000000000000"
   ,210 => "000000000000000000"
   ,211 => "000000000000000000"
   ,212 => "000000000000000000"
   ,213 => "000000000000000000"
   ,214 => "000000000000000000"
   ,215 => "000000000000000000"
   ,216 => "000000000000000000"
   ,217 => "000000000000000000"
   ,218 => "000000000000000000"
   ,219 => "000000000000000000"
   ,220 => "000000000000000000"
   ,221 => "000000000000000000"
   ,222 => "000000000000000000"
   ,223 => "000000000000000000"
   ,224 => "000000000000000000"
   ,225 => "000000000000000000"
   ,226 => "000000000000000000"
   ,227 => "000000000000000000"
   ,228 => "000000000000000000"
   ,229 => "000000000000000000"
   ,230 => "000000000000000000"
   ,231 => "000000000000000000"
   ,232 => "000000000000000000"
   ,233 => "000000000000000000"
   ,234 => "000000000000000000"
   ,235 => "000000000000000000"
   ,236 => "000000000000000000"
   ,237 => "000000000000000000"
   ,238 => "000000000000000000"
   ,239 => "000000000000000000"
   ,240 => "000000000000000000"
   ,241 => "000000000000000000"
   ,242 => "000000000000000000"
   ,243 => "000000000000000000"
   ,244 => "000000000000000000"
   ,245 => "000000000000000000"
   ,246 => "000000000000000000"
   ,247 => "000000000000000000"
   ,248 => "000000000000000000"
   ,249 => "000000000000000000"
   ,250 => "000000000000000000"
   ,251 => "000000000000000000"
   ,252 => "000000000000000000"
   ,253 => "000000000000000000"
   ,254 => "000000000000000000"
   ,255 => "000000000000000000"
   ,256 => "000000000000000000"
   ,257 => "000000000000000000"
   ,258 => "000000000000000000"
   ,259 => "000000000000000000"
   ,260 => "000000000000000000"
   ,261 => "000000000000000000"
   ,262 => "000000000000000000"
   ,263 => "000000000000000000"
   ,264 => "000000000000000000"
   ,265 => "000000000000000000"
   ,266 => "000000000000000000"
   ,267 => "000000000000000000"
   ,268 => "000000000000000000"
   ,269 => "000000000000000000"
   ,270 => "000000000000000000"
   ,271 => "000000000000000000"
   ,272 => "000000000000000000"
   ,273 => "000000000000000000"
   ,274 => "000000000000000000"
   ,275 => "000000000000000000"
   ,276 => "000000000000000000"
   ,277 => "000000000000000000"
   ,278 => "000000000000000000"
   ,279 => "000000000000000000"
   ,280 => "000000000000000000"
   ,281 => "000000000000000000"
   ,282 => "000000000000000000"
   ,283 => "000000000000000000"
   ,284 => "000000000000000000"
   ,285 => "000000000000000000"
   ,286 => "000000000000000000"
   ,287 => "000000000000000000"
   ,288 => "000000000000000000"
   ,289 => "000000000000000000"
   ,290 => "000000000000000000"
   ,291 => "000000000000000000"
   ,292 => "000000000000000000"
   ,293 => "000000000000000000"
   ,294 => "000000000000000000"
   ,295 => "000000000000000000"
   ,296 => "000000000000000000"
   ,297 => "000000000000000000"
   ,298 => "000000000000000000"
   ,299 => "000000000000000000"
   ,300 => "000000000000000000"
   ,301 => "000000000000000000"
   ,302 => "000000000000000000"
   ,303 => "000000000000000000"
   ,304 => "000000000000000000"
   ,305 => "000000000000000000"
   ,306 => "000000000000000000"
   ,307 => "000000000000000000"
   ,308 => "000000000000000000"
   ,309 => "000000000000000000"
   ,310 => "000000000000000000"
   ,311 => "000000000000000000"
   ,312 => "000000000000000000"
   ,313 => "000000000000000000"
   ,314 => "000000000000000000"
   ,315 => "000000000000000000"
   ,316 => "000000000000000000"
   ,317 => "000000000000000000"
   ,318 => "000000000000000000"
   ,319 => "000000000000000000"
   ,320 => "000000000000000000"
   ,321 => "000000000000000000"
   ,322 => "000000000000000000"
   ,323 => "000000000000000000"
   ,324 => "000000000000000000"
   ,325 => "000000000000000000"
   ,326 => "000000000000000000"
   ,327 => "000000000000000000"
   ,328 => "000000000000000000"
   ,329 => "000000000000000000"
   ,330 => "000000000000000000"
   ,331 => "000000000000000000"
   ,332 => "000000000000000000"
   ,333 => "000000000000000000"
   ,334 => "000000000000000000"
   ,335 => "000000000000000000"
   ,336 => "000000000000000000"
   ,337 => "000000000000000000"
   ,338 => "000000000000000000"
   ,339 => "000000000000000000"
   ,340 => "000000000000000000"
   ,341 => "000000000000000000"
   ,342 => "000000000000000000"
   ,343 => "000000000000000000"
   ,344 => "000000000000000000"
   ,345 => "000000000000000000"
   ,346 => "000000000000000000"
   ,347 => "000000000000000000"
   ,348 => "000000000000000000"
   ,349 => "000000000000000000"
   ,350 => "000000000000000000"
   ,351 => "000000000000000000"
   ,352 => "000000000000000000"
   ,353 => "000000000000000000"
   ,354 => "000000000000000000"
   ,355 => "000000000000000000"
   ,356 => "000000000000000000"
   ,357 => "000000000000000000"
   ,358 => "000000000000000000"
   ,359 => "000000000000000000"
   ,360 => "000000000000000000"
   ,361 => "000000000000000000"
   ,362 => "000000000000000000"
   ,363 => "000000000000000000"
   ,364 => "000000000000000000"
   ,365 => "000000000000000000"
   ,366 => "000000000000000000"
   ,367 => "000000000000000000"
   ,368 => "000000000000000000"
   ,369 => "000000000000000000"
   ,370 => "000000000000000000"
   ,371 => "000000000000000000"
   ,372 => "000000000000000000"
   ,373 => "000000000000000000"
   ,374 => "000000000000000000"
   ,375 => "000000000000000000"
   ,376 => "000000000000000000"
   ,377 => "000000000000000000"
   ,378 => "000000000000000000"
   ,379 => "000000000000000000"
   ,380 => "000000000000000000"
   ,381 => "000000000000000000"
   ,382 => "000000000000000000"
   ,383 => "000000000000000000"
   ,384 => "000000000000000000"
   ,385 => "000000000000000000"
   ,386 => "000000000000000000"
   ,387 => "000000000000000000"
   ,388 => "000000000000000000"
   ,389 => "000000000000000000"
   ,390 => "000000000000000000"
   ,391 => "000000000000000000"
   ,392 => "000000000000000000"
   ,393 => "000000000000000000"
   ,394 => "000000000000000000"
   ,395 => "000000000000000000"
   ,396 => "000000000000000000"
   ,397 => "000000000000000000"
   ,398 => "000000000000000000"
   ,399 => "000000000000000000"
   ,400 => "000000000000000000"
   ,401 => "000000000000000000"
   ,402 => "000000000000000000"
   ,403 => "000000000000000000"
   ,404 => "000000000000000000"
   ,405 => "000000000000000000"
   ,406 => "000000000000000000"
   ,407 => "000000000000000000"
   ,408 => "000000000000000000"
   ,409 => "000000000000000000"
   ,410 => "000000000000000000"
   ,411 => "000000000000000000"
   ,412 => "000000000000000000"
   ,413 => "000000000000000000"
   ,414 => "000000000000000000"
   ,415 => "000000000000000000"
   ,416 => "000000000000000000"
   ,417 => "000000000000000000"
   ,418 => "000000000000000000"
   ,419 => "000000000000000000"
   ,420 => "000000000000000000"
   ,421 => "000000000000000000"
   ,422 => "000000000000000000"
   ,423 => "000000000000000000"
   ,424 => "000000000000000000"
   ,425 => "000000000000000000"
   ,426 => "000000000000000000"
   ,427 => "000000000000000000"
   ,428 => "000000000000000000"
   ,429 => "000000000000000000"
   ,430 => "000000000000000000"
   ,431 => "000000000000000000"
   ,432 => "000000000000000000"
   ,433 => "000000000000000000"
   ,434 => "000000000000000000"
   ,435 => "000000000000000000"
   ,436 => "000000000000000000"
   ,437 => "000000000000000000"
   ,438 => "000000000000000000"
   ,439 => "000000000000000000"
   ,440 => "000000000000000000"
   ,441 => "000000000000000000"
   ,442 => "000000000000000000"
   ,443 => "000000000000000000"
   ,444 => "000000000000000000"
   ,445 => "000000000000000000"
   ,446 => "000000000000000000"
   ,447 => "000000000000000000"
   ,448 => "000000000000000000"
   ,449 => "000000000000000000"
   ,450 => "000000000000000000"
   ,451 => "000000000000000000"
   ,452 => "000000000000000000"
   ,453 => "000000000000000000"
   ,454 => "000000000000000000"
   ,455 => "000000000000000000"
   ,456 => "000000000000000000"
   ,457 => "000000000000000000"
   ,458 => "000000000000000000"
   ,459 => "000000000000000000"
   ,460 => "000000000000000000"
   ,461 => "000000000000000000"
   ,462 => "000000000000000000"
   ,463 => "000000000000000000"
   ,464 => "000000000000000000"
   ,465 => "000000000000000000"
   ,466 => "000000000000000000"
   ,467 => "000000000000000000"
   ,468 => "000000000000000000"
   ,469 => "000000000000000000"
   ,470 => "000000000000000000"
   ,471 => "000000000000000000"
   ,472 => "000000000000000000"
   ,473 => "000000000000000000"
   ,474 => "000000000000000000"
   ,475 => "000000000000000000"
   ,476 => "000000000000000000"
   ,477 => "000000000000000000"
   ,478 => "000000000000000000"
   ,479 => "000000000000000000"
   ,480 => "000000000000000000"
   ,481 => "000000000000000000"
   ,482 => "000000000000000000"
   ,483 => "000000000000000000"
   ,484 => "000000000000000000"
   ,485 => "000000000000000000"
   ,486 => "000000000000000000"
   ,487 => "000000000000000000"
   ,488 => "000000000000000000"
   ,489 => "000000000000000000"
   ,490 => "000000000000000000"
   ,491 => "000000000000000000"
   ,492 => "000000000000000000"
   ,493 => "000000000000000000"
   ,494 => "000000000000000000"
   ,495 => "000000000000000000"
   ,496 => "000000000000000000"
   ,497 => "000000000000000000"
   ,498 => "000000000000000000"
   ,499 => "000000000000000000"
   ,500 => "000000000000000000"
   ,501 => "000000000000000000"
   ,502 => "000000000000000000"
   ,503 => "000000000000000000"
   ,504 => "000000000000000000"
   ,505 => "000000000000000000"
   ,506 => "000000000000000000"
   ,507 => "000000000000000000"
   ,508 => "000000000000000000"
   ,509 => "000000000000000000"
   ,510 => "000000000000000000"
   ,511 => "000000000000000000"
   ,512 => "000000000000000000"
   ,513 => "000000000000000000"
   ,514 => "000000000000000000"
   ,515 => "000000000000000000"
   ,516 => "000000000000000000"
   ,517 => "000000000000000000"
   ,518 => "000000000000000000"
   ,519 => "000000000000000000"
   ,520 => "000000000000000000"
   ,521 => "000000000000000000"
   ,522 => "000000000000000000"
   ,523 => "000000000000000000"
   ,524 => "000000000000000000"
   ,525 => "000000000000000000"
   ,526 => "000000000000000000"
   ,527 => "000000000000000000"
   ,528 => "000000000000000000"
   ,529 => "000000000000000000"
   ,530 => "000000000000000000"
   ,531 => "000000000000000000"
   ,532 => "000000000000000000"
   ,533 => "000000000000000000"
   ,534 => "000000000000000000"
   ,535 => "000000000000000000"
   ,536 => "000000000000000000"
   ,537 => "000000000000000000"
   ,538 => "000000000000000000"
   ,539 => "000000000000000000"
   ,540 => "000000000000000000"
   ,541 => "000000000000000000"
   ,542 => "000000000000000000"
   ,543 => "000000000000000000"
   ,544 => "000000000000000000"
   ,545 => "000000000000000000"
   ,546 => "000000000000000000"
   ,547 => "000000000000000000"
   ,548 => "000000000000000000"
   ,549 => "000000000000000000"
   ,550 => "000000000000000000"
   ,551 => "000000000000000000"
   ,552 => "000000000000000000"
   ,553 => "000000000000000000"
   ,554 => "000000000000000000"
   ,555 => "000000000000000000"
   ,556 => "000000000000000000"
   ,557 => "000000000000000000"
   ,558 => "000000000000000000"
   ,559 => "000000000000000000"
   ,560 => "000000000000000000"
   ,561 => "000000000000000000"
   ,562 => "000000000000000000"
   ,563 => "000000000000000000"
   ,564 => "000000000000000000"
   ,565 => "000000000000000000"
   ,566 => "000000000000000000"
   ,567 => "000000000000000000"
   ,568 => "000000000000000000"
   ,569 => "000000000000000000"
   ,570 => "000000000000000000"
   ,571 => "000000000000000000"
   ,572 => "000000000000000000"
   ,573 => "000000000000000000"
   ,574 => "000000000000000000"
   ,575 => "000000000000000000"
   ,576 => "000000000000000000"
   ,577 => "000000000000000000"
   ,578 => "000000000000000000"
   ,579 => "000000000000000000"
   ,580 => "000000000000000000"
   ,581 => "000000000000000000"
   ,582 => "000000000000000000"
   ,583 => "000000000000000000"
   ,584 => "000000000000000000"
   ,585 => "000000000000000000"
   ,586 => "000000000000000000"
   ,587 => "000000000000000000"
   ,588 => "000000000000000000"
   ,589 => "000000000000000000"
   ,590 => "000000000000000000"
   ,591 => "000000000000000000"
   ,592 => "000000000000000000"
   ,593 => "000000000000000000"
   ,594 => "000000000000000000"
   ,595 => "000000000000000000"
   ,596 => "000000000000000000"
   ,597 => "000000000000000000"
   ,598 => "000000000000000000"
   ,599 => "000000000000000000"
   ,600 => "000000000000000000"
   ,601 => "000000000000000000"
   ,602 => "000000000000000000"
   ,603 => "000000000000000000"
   ,604 => "000000000000000000"
   ,605 => "000000000000000000"
   ,606 => "000000000000000000"
   ,607 => "000000000000000000"
   ,608 => "000000000000000000"
   ,609 => "000000000000000000"
   ,610 => "000000000000000000"
   ,611 => "000000000000000000"
   ,612 => "000000000000000000"
   ,613 => "000000000000000000"
   ,614 => "000000000000000000"
   ,615 => "000000000000000000"
   ,616 => "000000000000000000"
   ,617 => "000000000000000000"
   ,618 => "000000000000000000"
   ,619 => "000000000000000000"
   ,620 => "000000000000000000"
   ,621 => "000000000000000000"
   ,622 => "000000000000000000"
   ,623 => "000000000000000000"
   ,624 => "000000000000000000"
   ,625 => "000000000000000000"
   ,626 => "000000000000000000"
   ,627 => "000000000000000000"
   ,628 => "000000000000000000"
   ,629 => "000000000000000000"
   ,630 => "000000000000000000"
   ,631 => "000000000000000000"
   ,632 => "000000000000000000"
   ,633 => "000000000000000000"
   ,634 => "000000000000000000"
   ,635 => "000000000000000000"
   ,636 => "000000000000000000"
   ,637 => "000000000000000000"
   ,638 => "000000000000000000"
   ,639 => "000000000000000000"
   ,640 => "000000000000000000"
   ,641 => "000000000000000000"
   ,642 => "000000000000000000"
   ,643 => "000000000000000000"
   ,644 => "000000000000000000"
   ,645 => "000000000000000000"
   ,646 => "000000000000000000"
   ,647 => "000000000000000000"
   ,648 => "000000000000000000"
   ,649 => "000000000000000000"
   ,650 => "000000000000000000"
   ,651 => "000000000000000000"
   ,652 => "000000000000000000"
   ,653 => "000000000000000000"
   ,654 => "000000000000000000"
   ,655 => "000000000000000000"
   ,656 => "000000000000000000"
   ,657 => "000000000000000000"
   ,658 => "000000000000000000"
   ,659 => "000000000000000000"
   ,660 => "000000000000000000"
   ,661 => "000000000000000000"
   ,662 => "000000000000000000"
   ,663 => "000000000000000000"
   ,664 => "000000000000000000"
   ,665 => "000000000000000000"
   ,666 => "000000000000000000"
   ,667 => "000000000000000000"
   ,668 => "000000000000000000"
   ,669 => "000000000000000000"
   ,670 => "000000000000000000"
   ,671 => "000000000000000000"
   ,672 => "000000000000000000"
   ,673 => "000000000000000000"
   ,674 => "000000000000000000"
   ,675 => "000000000000000000"
   ,676 => "000000000000000000"
   ,677 => "000000000000000000"
   ,678 => "000000000000000000"
   ,679 => "000000000000000000"
   ,680 => "000000000000000000"
   ,681 => "000000000000000000"
   ,682 => "000000000000000000"
   ,683 => "000000000000000000"
   ,684 => "000000000000000000"
   ,685 => "000000000000000000"
   ,686 => "000000000000000000"
   ,687 => "000000000000000000"
   ,688 => "000000000000000000"
   ,689 => "000000000000000000"
   ,690 => "000000000000000000"
   ,691 => "000000000000000000"
   ,692 => "000000000000000000"
   ,693 => "000000000000000000"
   ,694 => "000000000000000000"
   ,695 => "000000000000000000"
   ,696 => "000000000000000000"
   ,697 => "000000000000000000"
   ,698 => "000000000000000000"
   ,699 => "000000000000000000"
   ,700 => "000000000000000000"
   ,701 => "000000000000000000"
   ,702 => "000000000000000000"
   ,703 => "000000000000000000"
   ,704 => "000000000000000000"
   ,705 => "000000000000000000"
   ,706 => "000000000000000000"
   ,707 => "000000000000000000"
   ,708 => "000000000000000000"
   ,709 => "000000000000000000"
   ,710 => "000000000000000000"
   ,711 => "000000000000000000"
   ,712 => "000000000000000000"
   ,713 => "000000000000000000"
   ,714 => "000000000000000000"
   ,715 => "000000000000000000"
   ,716 => "000000000000000000"
   ,717 => "000000000000000000"
   ,718 => "000000000000000000"
   ,719 => "000000000000000000"
   ,720 => "000000000000000000"
   ,721 => "000000000000000000"
   ,722 => "000000000000000000"
   ,723 => "000000000000000000"
   ,724 => "000000000000000000"
   ,725 => "000000000000000000"
   ,726 => "000000000000000000"
   ,727 => "000000000000000000"
   ,728 => "000000000000000000"
   ,729 => "000000000000000000"
   ,730 => "000000000000000000"
   ,731 => "000000000000000000"
   ,732 => "000000000000000000"
   ,733 => "000000000000000000"
   ,734 => "000000000000000000"
   ,735 => "000000000000000000"
   ,736 => "000000000000000000"
   ,737 => "000000000000000000"
   ,738 => "000000000000000000"
   ,739 => "000000000000000000"
   ,740 => "000000000000000000"
   ,741 => "000000000000000000"
   ,742 => "000000000000000000"
   ,743 => "000000000000000000"
   ,744 => "000000000000000000"
   ,745 => "000000000000000000"
   ,746 => "000000000000000000"
   ,747 => "000000000000000000"
   ,748 => "000000000000000000"
   ,749 => "000000000000000000"
   ,750 => "000000000000000000"
   ,751 => "000000000000000000"
   ,752 => "000000000000000000"
   ,753 => "000000000000000000"
   ,754 => "000000000000000000"
   ,755 => "000000000000000000"
   ,756 => "000000000000000000"
   ,757 => "000000000000000000"
   ,758 => "000000000000000000"
   ,759 => "000000000000000000"
   ,760 => "000000000000000000"
   ,761 => "000000000000000000"
   ,762 => "000000000000000000"
   ,763 => "000000000000000000"
   ,764 => "000000000000000000"
   ,765 => "000000000000000000"
   ,766 => "000000000000000000"
   ,767 => "000000000000000000"
   ,768 => "000000000000000000"
   ,769 => "000000000000000000"
   ,770 => "000000000000000000"
   ,771 => "000000000000000000"
   ,772 => "000000000000000000"
   ,773 => "000000000000000000"
   ,774 => "000000000000000000"
   ,775 => "000000000000000000"
   ,776 => "000000000000000000"
   ,777 => "000000000000000000"
   ,778 => "000000000000000000"
   ,779 => "000000000000000000"
   ,780 => "000000000000000000"
   ,781 => "000000000000000000"
   ,782 => "000000000000000000"
   ,783 => "000000000000000000"
   ,784 => "000000000000000000"
   ,785 => "000000000000000000"
   ,786 => "000000000000000000"
   ,787 => "000000000000000000"
   ,788 => "000000000000000000"
   ,789 => "000000000000000000"
   ,790 => "000000000000000000"
   ,791 => "000000000000000000"
   ,792 => "000000000000000000"
   ,793 => "000000000000000000"
   ,794 => "000000000000000000"
   ,795 => "000000000000000000"
   ,796 => "000000000000000000"
   ,797 => "000000000000000000"
   ,798 => "000000000000000000"
   ,799 => "000000000000000000"
   ,800 => "000000000000000000"
   ,801 => "000000000000000000"
   ,802 => "000000000000000000"
   ,803 => "000000000000000000"
   ,804 => "000000000000000000"
   ,805 => "000000000000000000"
   ,806 => "000000000000000000"
   ,807 => "000000000000000000"
   ,808 => "000000000000000000"
   ,809 => "000000000000000000"
   ,810 => "000000000000000000"
   ,811 => "000000000000000000"
   ,812 => "000000000000000000"
   ,813 => "000000000000000000"
   ,814 => "000000000000000000"
   ,815 => "000000000000000000"
   ,816 => "000000000000000000"
   ,817 => "000000000000000000"
   ,818 => "000000000000000000"
   ,819 => "000000000000000000"
   ,820 => "000000000000000000"
   ,821 => "000000000000000000"
   ,822 => "000000000000000000"
   ,823 => "000000000000000000"
   ,824 => "000000000000000000"
   ,825 => "000000000000000000"
   ,826 => "000000000000000000"
   ,827 => "000000000000000000"
   ,828 => "000000000000000000"
   ,829 => "000000000000000000"
   ,830 => "000000000000000000"
   ,831 => "000000000000000000"
   ,832 => "000000000000000000"
   ,833 => "000000000000000000"
   ,834 => "000000000000000000"
   ,835 => "000000000000000000"
   ,836 => "000000000000000000"
   ,837 => "000000000000000000"
   ,838 => "000000000000000000"
   ,839 => "000000000000000000"
   ,840 => "000000000000000000"
   ,841 => "000000000000000000"
   ,842 => "000000000000000000"
   ,843 => "000000000000000000"
   ,844 => "000000000000000000"
   ,845 => "000000000000000000"
   ,846 => "000000000000000000"
   ,847 => "000000000000000000"
   ,848 => "000000000000000000"
   ,849 => "000000000000000000"
   ,850 => "000000000000000000"
   ,851 => "000000000000000000"
   ,852 => "000000000000000000"
   ,853 => "000000000000000000"
   ,854 => "000000000000000000"
   ,855 => "000000000000000000"
   ,856 => "000000000000000000"
   ,857 => "000000000000000000"
   ,858 => "000000000000000000"
   ,859 => "000000000000000000"
   ,860 => "000000000000000000"
   ,861 => "000000000000000000"
   ,862 => "000000000000000000"
   ,863 => "000000000000000000"
   ,864 => "000000000000000000"
   ,865 => "000000000000000000"
   ,866 => "000000000000000000"
   ,867 => "000000000000000000"
   ,868 => "000000000000000000"
   ,869 => "000000000000000000"
   ,870 => "000000000000000000"
   ,871 => "000000000000000000"
   ,872 => "000000000000000000"
   ,873 => "000000000000000000"
   ,874 => "000000000000000000"
   ,875 => "000000000000000000"
   ,876 => "000000000000000000"
   ,877 => "000000000000000000"
   ,878 => "000000000000000000"
   ,879 => "000000000000000000"
   ,880 => "000000000000000000"
   ,881 => "000000000000000000"
   ,882 => "000000000000000000"
   ,883 => "000000000000000000"
   ,884 => "000000000000000000"
   ,885 => "000000000000000000"
   ,886 => "000000000000000000"
   ,887 => "000000000000000000"
   ,888 => "000000000000000000"
   ,889 => "000000000000000000"
   ,890 => "000000000000000000"
   ,891 => "000000000000000000"
   ,892 => "000000000000000000"
   ,893 => "000000000000000000"
   ,894 => "000000000000000000"
   ,895 => "000000000000000000"
   ,896 => "000000000000000000"
   ,897 => "000000000000000000"
   ,898 => "000000000000000000"
   ,899 => "000000000000000000"
   ,900 => "000000000000000000"
   ,901 => "000000000000000000"
   ,902 => "000000000000000000"
   ,903 => "000000000000000000"
   ,904 => "000000000000000000"
   ,905 => "000000000000000000"
   ,906 => "000000000000000000"
   ,907 => "000000000000000000"
   ,908 => "000000000000000000"
   ,909 => "000000000000000000"
   ,910 => "000000000000000000"
   ,911 => "000000000000000000"
   ,912 => "000000000000000000"
   ,913 => "000000000000000000"
   ,914 => "000000000000000000"
   ,915 => "000000000000000000"
   ,916 => "000000000000000000"
   ,917 => "000000000000000000"
   ,918 => "000000000000000000"
   ,919 => "000000000000000000"
   ,920 => "000000000000000000"
   ,921 => "000000000000000000"
   ,922 => "000000000000000000"
   ,923 => "000000000000000000"
   ,924 => "000000000000000000"
   ,925 => "000000000000000000"
   ,926 => "000000000000000000"
   ,927 => "000000000000000000"
   ,928 => "000000000000000000"
   ,929 => "000000000000000000"
   ,930 => "000000000000000000"
   ,931 => "000000000000000000"
   ,932 => "000000000000000000"
   ,933 => "000000000000000000"
   ,934 => "000000000000000000"
   ,935 => "000000000000000000"
   ,936 => "000000000000000000"
   ,937 => "000000000000000000"
   ,938 => "000000000000000000"
   ,939 => "000000000000000000"
   ,940 => "000000000000000000"
   ,941 => "000000000000000000"
   ,942 => "000000000000000000"
   ,943 => "000000000000000000"
   ,944 => "000000000000000000"
   ,945 => "000000000000000000"
   ,946 => "000000000000000000"
   ,947 => "000000000000000000"
   ,948 => "000000000000000000"
   ,949 => "000000000000000000"
   ,950 => "000000000000000000"
   ,951 => "000000000000000000"
   ,952 => "000000000000000000"
   ,953 => "000000000000000000"
   ,954 => "000000000000000000"
   ,955 => "000000000000000000"
   ,956 => "000000000000000000"
   ,957 => "000000000000000000"
   ,958 => "000000000000000000"
   ,959 => "000000000000000000"
   ,960 => "000000000000000000"
   ,961 => "000000000000000000"
   ,962 => "000000000000000000"
   ,963 => "000000000000000000"
   ,964 => "000000000000000000"
   ,965 => "000000000000000000"
   ,966 => "000000000000000000"
   ,967 => "000000000000000000"
   ,968 => "000000000000000000"
   ,969 => "000000000000000000"
   ,970 => "000000000000000000"
   ,971 => "000000000000000000"
   ,972 => "000000000000000000"
   ,973 => "000000000000000000"
   ,974 => "000000000000000000"
   ,975 => "000000000000000000"
   ,976 => "000000000000000000"
   ,977 => "000000000000000000"
   ,978 => "000000000000000000"
   ,979 => "000000000000000000"
   ,980 => "000000000000000000"
   ,981 => "000000000000000000"
   ,982 => "000000000000000000"
   ,983 => "000000000000000000"
   ,984 => "000000000000000000"
   ,985 => "000000000000000000"
   ,986 => "000000000000000000"
   ,987 => "000000000000000000"
   ,988 => "000000000000000000"
   ,989 => "000000000000000000"
   ,990 => "000000000000000000"
   ,991 => "000000000000000000"
   ,992 => "000000000000000000"
   ,993 => "000000000000000000"
   ,994 => "000000000000000000"
   ,995 => "000000000000000000"
   ,996 => "000000000000000000"
   ,997 => "000000000000000000"
   ,998 => "000000000000000000"
   ,999 => "000000000000000000"
   ,1000 => "000000000000000000"
   ,1001 => "000000000000000000"
   ,1002 => "000000000000000000"
   ,1003 => "000000000000000000"
   ,1004 => "000000000000000000"
   ,1005 => "000000000000000000"
   ,1006 => "000000000000000000"
   ,1007 => "000000000000000000"
   ,1008 => "000000000000000000"
   ,1009 => "000000000000000000"
   ,1010 => "000000000000000000"
   ,1011 => "000000000000000000"
   ,1012 => "000000000000000000"
   ,1013 => "000000000000000000"
   ,1014 => "000000000000000000"
   ,1015 => "000000000000000000"
   ,1016 => "000000000000000000"
   ,1017 => "000000000000000000"
   ,1018 => "000000000000000000"
   ,1019 => "000000000000000000"
   ,1020 => "000000000000000000"
   ,1021 => "000000000000000000"
   ,1022 => "000000000000000000"
   ,1023 => "111000000000000001"
   );
begin
  process(clk_i)
  begin
    if(clk_i'event and clk_i = '1') then
       data_o <= rom(to_integer(unsigned(addr_i)));
    end if;
  end process;
end rtl;
