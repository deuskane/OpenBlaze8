-------------------------------------------------------------------------------
-- Title      : vga_font_memory
-- Project    : PicoSOC
-------------------------------------------------------------------------------
-- File       : vga_font_memory.vhd
-- Author     : Mathieu Rosière
-- Company    : 
-- Created    : 2014-01-04
-- Last update: 2017-03-31
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2013 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-01-04  0.1      rosière	Created
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity vga_font_memory is
  generic(DEPTH_MAX      : natural := 2**8;  -- ASCII : 8bits
          SIZE_CHAR_X_MAX: natural := 8;
          SIZE_CHAR_Y_MAX: natural := 16;
          SIZE_ADDR_ID   : natural := 8;
          SIZE_ADDR_X    : natural := 3;
          SIZE_ADDR_Y    : natural := 4
          );
  port   (
--        clk_i          : in   std_logic;
--        arstn_i        : in   std_logic;

          character_id_i : in   std_logic_vector(SIZE_ADDR_ID-1 downto 0);
          character_x_i  : in   std_logic_vector(SIZE_ADDR_X-1  downto 0);
          character_y_i  : in   std_logic_vector(SIZE_ADDR_Y-1  downto 0);
          
          pixel_o        : out  std_logic
          );
end vga_font_memory;

architecture rtl of vga_font_memory is
  -- =====[ Types ]===============================
  type character_t    is array (0 to SIZE_CHAR_Y_MAX-1) of std_logic_vector(0 to SIZE_CHAR_X_MAX-1);
  type font_memory_t  is array (DEPTH_MAX-1 downto 0) of character_t;

  -- =====[ Registers ]===========================
  
  -- =====[ Signals ]=============================
  --signal   font_memory_r           : font_memory_t;
  constant font_memory_r           : font_memory_t :=
    --         x: 0      7
    (-- d000 - x00 - NUL
     0       => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d037 - x25 - '%'
    , 37     => ("00000000" -- y=0
                ,"00000000"
                ,"01100110"
                ,"01100110"
                ,"00001100"
                ,"00001100"
                ,"00001000"
                ,"00011000"
                ,"00011000"
                ,"00010000"
                ,"00110000"
                ,"00110000"
                ,"01100110"
                ,"01100110"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d042 - x2a - '*'
    , 42     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00011000"
                ,"00011000"
                ,"01111110"
                ,"00111100"
                ,"00011000"
                ,"00100100"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d043 - x2b - '+'
    , 43     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00011000"
                ,"00011000"
                ,"01111110"
                ,"01111110"
                ,"00011000"
                ,"00011000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d045 - x2d - '-'
    , 45     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d047 - x2f - '/'
    , 47     => ("00000000" -- y=0
                ,"00000000"
                ,"00000110"
                ,"00000110"
                ,"00001100"
                ,"00001100"
                ,"00001000"
                ,"00011000"
                ,"00011000"
                ,"00010000"
                ,"00110000"
                ,"00110000"
                ,"01100000"
                ,"01100000"
                ,"00000000"
                ,"00000000" -- y=15
                 )


     
    -- d048 - x30 - '0'
    , 48     => ("00000000" -- y=0
                ,"00000000"
                ,"00111100"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"00111100"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d049 - x31 - '1'
    , 49     => ("00000000" -- y=0
                ,"00000000"
                ,"00011000"
                ,"00111000"
                ,"01111000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d050 - x32 - '2'
    , 50     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"01111110"
                ,"01111110"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d051 - x33 - '3'
    , 51     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"00011110"
                ,"00011110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d052 - x34 - '4'
    , 52     => ("00000000" -- y=0
                ,"00000000"
                ,"00001100"
                ,"00011100"
                ,"00111100"
                ,"00101100"
                ,"00101100"
                ,"01101100"
                ,"01101100"
                ,"01111110"
                ,"01111110"
                ,"00001100"
                ,"00001100"
                ,"00001100"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d053 - x35 - '5'
    , 53     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01111110"
                ,"01111110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d054 - x36 - '6'
    , 54     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01111110"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d055 - x37 - '7'
    , 55     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"00000110"
                ,"00000110"
                ,"00001100"
                ,"00001100"
                ,"00011000"
                ,"00011000"
                ,"00110000"
                ,"00110000"
                ,"01100000"
                ,"01100000"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d056 - x38 - '8'
    , 56     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d057 - x39 - '9'
    , 57     => ("00000000" -- y=0
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"01111110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d061 - x3D - '='
    , 61     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000"
                ,"01111110"
                ,"01111110"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000" -- y=15
                 )

    -- d097 - x61 - 'a'
    , 97     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"01111100"
                ,"01111110"
                ,"00000110"
                ,"00000110"
                ,"00111110"
                ,"01100110"
                ,"01111110"
                ,"00111010"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d098 - x62 - 'b'
    , 98     => ("00000000" -- y=0
                ,"00000000"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01111100"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"01111100"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d099 - x63 - 'c'
    , 99     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00111110"
                ,"01111110"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01100000"
                ,"01111110"
                ,"00111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d100 - x64 - 'd'
    ,100     => ("00000000" -- y=0
                ,"00000000"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"00000110"
                ,"00111110"
                ,"01111110"
                ,"01100110"
                ,"01100110"
                ,"01111110"
                ,"00111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d101 - x65 - 'e'
    ,101     => ("00000000" -- y=0
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00000000"
                ,"00111100"
                ,"01111110"
                ,"01100110"
                ,"01111110"
                ,"01100000"
                ,"01100000"
                ,"01111110"
                ,"00111110"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- d102 - x66 - 'f'
    ,102     => ("00000000" -- y=0
                ,"00000000"
                ,"00001110"
                ,"00011110"
                ,"00011000"
                ,"00011000"
                ,"01111110"
                ,"01111110"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00000000"
                ,"00000000" -- y=15
                 )
     
    -- others : X
    ,others  => ("10000001" -- y=0
                ,"10000001"
                ,"01000010"
                ,"01000010"
                ,"00100100"
                ,"00100100"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00011000"
                ,"00100100"
                ,"00100100"
                ,"01000010"
                ,"01000010"
                ,"10000001"
                ,"10000001" -- y=15
                 )

     );

begin


  pixel_o <= font_memory_r(to_integer(unsigned(character_id_i)))
                          (to_integer(unsigned(character_y_i )))
                          (to_integer(unsigned(character_x_i )));
  
end rtl;
